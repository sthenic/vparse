reg a_register;
