module A();

    B B_inst ();
    C C_inst ();

endmodule
