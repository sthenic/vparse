module modB();

    modD();
    modC();

endmodule
