module B();

    D D_inst ();
    E E_inst ();

endmodule
