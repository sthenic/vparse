module G();
endmodule
