wire wire2;
`include "test3.vh"
wire next_to_last_wire;
