`define WIDTH 8
