`__FILE__
