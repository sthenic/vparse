wire wire3;
