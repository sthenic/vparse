module modD();

endmodule
