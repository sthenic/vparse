


`__LINE__
