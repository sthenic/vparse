module needs_includemod();

    includemod includemod_inst();

endmodule
