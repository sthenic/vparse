module C();
endmodule
