module modA();

    modC();
    modD();
    modB();

endmodule
