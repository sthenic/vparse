module modC();

    modD();

endmodule
