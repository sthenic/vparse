wire [7:0] my_wire;
