module includemod();

endmodule
