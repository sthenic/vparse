module H();

endmodule
