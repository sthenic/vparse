module D();
endmodule

module E();
endmodule
