module F();

    G G_inst ();
    B B_inst ();

endmodule
