`FOO my_reg;
